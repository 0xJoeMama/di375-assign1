library ieee;
use ieee.std_logic_1164.all;


entity majority is
  port(
  a, b, c: in STD_LOGIC;
  y: out STD_LOGIC
  );
end entity majority;

architecture dataflow of majority is
begin
  y <= (a and (b or c)) or (b and c);
end architecture dataflow;
